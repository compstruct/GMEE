
module Mult4(product,inp1,inp2);
output [7:0]product;
input [3:0]inp1;
input [3:0]inp2;
assign product[0]=(inp1[0]&inp2[0]);
wire x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,x16,x17;

HA1 HA1(product[1],x1,(inp1[1]&inp2[0]),(inp1[0]&inp2[1]));
FA1 FA1(x2,x3,inp1[1]&inp2[1],(inp1[0]&inp2[2]),x1);
FA1 FA2(x4,x5,(inp1[1]&inp2[2]),(inp1[0]&inp2[3]),x3);
HA1 HA2(x6,x7,(inp1[1]&inp2[3]),x5);

HA1 HA3(product[2],x15,x2,(inp1[2]&inp2[0]));
FA1 FA5(x14,x16,x4,(inp1[2]&inp2[1]),x15);
FA1 FA4(x13,x17,x6,(inp1[2]&inp2[2]),x16);
FA1 FA3(x9,x8,x7,(inp1[2]&inp2[3]),x17);

HA1 HA4(product[3],x12,x14,(inp1[3]&inp2[0]));
FA1 FA8(product[4],x11,x13,(inp1[3]&inp2[1]),x12);
FA1 FA7(product[5],x10,x9,(inp1[3]&inp2[2]),x11);
FA1 FA6(product[6],product[7],x8,(inp1[3]&inp2[3]),x10);

endmodule



module Mult4_TT3(product,inp1,inp2); //replace the last line with TT3 FA
output [7:0]product;
input [3:0]inp1;
input [3:0]inp2;
assign product[0]=(inp1[0]&inp2[0]);
wire x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,x16,x17;
wire [7:0] accurate_product;

HA1_TT3 HA1(product[1],x1,(inp1[1]&inp2[0]),(inp1[0]&inp2[1]));
FA1_TT3 FA1(x2,x3,inp1[1]&inp2[1],(inp1[0]&inp2[2]),x1);
FA1_TT3 FA2(x4,x5,(inp1[1]&inp2[2]),(inp1[0]&inp2[3]),x3);
HA1 HA2(x6,x7,(inp1[1]&inp2[3]),x5);

HA1_TT3 HA3(product[2],x15,x2,(inp1[2]&inp2[0]));
FA1_TT3 FA5(x14,x16,x4,(inp1[2]&inp2[1]),x15);
FA1 FA4(x13,x17,x6,(inp1[2]&inp2[2]),x16);
FA1 FA3(x9,x8,x7,(inp1[2]&inp2[3]),x17);

HA1_TT3 HA4(product[3],x12,x14,(inp1[3]&inp2[0]));
FA1 FA8(product[4],x11,x13,(inp1[3]&inp2[1]),x12);
FA1 FA7(product[5],x10,x9,(inp1[3]&inp2[2]),x11);
FA1 FA6(product[6],product[7],x8,(inp1[3]&inp2[3]),x10);


//
assign accurate_product = inp1*inp2;
//


endmodule